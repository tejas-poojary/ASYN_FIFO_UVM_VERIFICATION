package async_fifo_pkg;
  import uvm_pkg::*;
 `include "uvm_macros.svh"
 `include "async_fifo_defines.sv"
 `include "async_fifo_wr_sequence_item.sv"
 `include "async_fifo_rd_sequence_item.sv"
 `include "async_fifo_wr_sequence.sv"
 `include "async_fifo_rd_sequence.sv"
 `include "async_fifo_wr_sequencer.sv"
 `include "async_fifo_rd_sequencer.sv"
 `include "async_fifo_wr_driver.sv"
 `include "async_fifo_rd_driver.sv"
 `include "async_fifo_wr_monitor.sv"
 `include "async_fifo_rd_monitor.sv"
 `include "async_fifo_wr_agent.sv"
 `include "async_fifo_rd_agent.sv"
 `include "async_fifo_subscriber.sv"
 `include "async_fifo_scoreboard.sv"
 `include "async_fifo_virtual_sequencer.sv"
 `include "async_fifo_virtual_sequence.sv"
 `include "async_fifo_environment.sv"
 `include "async_fifo_test.sv"
endpackage
