`define no_of_times 20
`define DSIZE 8
`define ASIZE 4
